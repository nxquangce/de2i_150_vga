module draw_superpixel();

endmodule